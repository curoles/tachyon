/* Writeback pipeline stage.
 *
 * Author:    Igor Lesik 2021
 * Copyright: Igor Lesik 2021
 *
 */
module Writeback #(
    parameter   ADDR_WIDTH = 32,
    localparam  ADDR_START = 2, // 4 bytes aligned
    localparam  INSN_SIZE  = 4,
    localparam  INSN_WIDTH = INSN_SIZE * 8
)(
    input  wire                           clk,
    input  wire                           rst,
    input  stage::InsnBundle              insn
);

    always @(posedge clk)
    begin
        if (!rst) begin
            $display("%4t WRB: addr=%h op=%h",
                $time, {insn.addr, 2'b00}, insn.insn);
        end else begin
            //
        end

    end


endmodule