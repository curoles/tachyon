`include "logmsg.svh"

/* Writeback pipeline stage.
 *
 * Author:    Igor Lesik 2021
 * Copyright: Igor Lesik 2021
 *
 */
module Writeback #(
    parameter   ADDR_WIDTH = stage::ADDR_WIDTH,
    localparam  ADDR_START = stage::ADDR_START,
    localparam  INSN_SIZE  = stage::INSN_SIZE,
    localparam  INSN_WIDTH = stage::INSN_WIDTH
)(
    input  wire                           clk,
    input  wire                           rst,
    input  stage::InsnBundle              insn
);

    always @(posedge clk)
    begin
        if (!rst) begin
            `MSG(5, ("WRB: addr=%h op=%h",
                {insn.addr, 2'b00}, insn.insn));
        end else begin
            //
        end

    end


endmodule